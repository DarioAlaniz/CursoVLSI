magic
tech sky130A
magscale 1 2
timestamp 1615311486
<< nwell >>
rect -525 517 -160 861
rect -525 485 -405 517
rect -374 485 -160 517
rect -525 484 -493 485
rect -366 484 -160 485
rect -525 476 -160 484
rect -525 475 -227 476
rect -220 475 -160 476
rect -525 470 -160 475
<< psubdiff >>
rect -480 -11 -456 23
rect -216 -11 -192 23
<< nsubdiff >>
rect -487 788 -463 822
rect -223 788 -199 822
<< psubdiffcont >>
rect -456 -11 -216 23
<< nsubdiffcont >>
rect -463 788 -223 822
<< poly >>
rect -405 375 -375 513
rect -470 364 -375 375
rect -470 330 -452 364
rect -418 330 -375 364
rect -470 318 -375 330
rect -405 295 -375 318
rect -317 449 -287 540
rect -317 438 -247 449
rect -317 404 -299 438
rect -265 404 -247 438
rect -317 392 -247 404
rect -317 284 -287 392
<< polycont >>
rect -452 330 -418 364
rect -299 404 -265 438
<< locali >>
rect -317 439 -248 448
rect -317 403 -300 439
rect -264 403 -248 439
rect -317 393 -248 403
rect -470 365 -401 374
rect -470 329 -453 365
rect -417 329 -401 365
rect -470 319 -401 329
<< viali >>
rect -487 788 -463 822
rect -463 788 -223 822
rect -223 788 -199 822
rect -300 438 -264 439
rect -300 404 -299 438
rect -299 404 -265 438
rect -265 404 -264 438
rect -300 403 -264 404
rect -453 364 -417 365
rect -453 330 -452 364
rect -452 330 -418 364
rect -418 330 -417 364
rect -453 329 -417 330
rect -480 -11 -456 23
rect -456 -11 -216 23
rect -216 -11 -192 23
<< metal1 >>
rect -525 822 -160 829
rect -525 788 -487 822
rect -199 788 -160 822
rect -525 782 -160 788
rect -454 550 -412 782
rect -360 570 -332 674
rect -361 505 -331 570
rect -276 550 -234 782
rect -361 477 -192 505
rect -227 476 -192 477
rect -317 439 -248 448
rect -317 431 -300 439
rect -525 403 -300 431
rect -264 403 -248 439
rect -317 393 -248 403
rect -470 365 -401 374
rect -470 357 -453 365
rect -525 329 -453 357
rect -417 329 -401 365
rect -220 332 -192 476
rect -470 321 -401 329
rect -272 303 -160 332
rect -451 29 -417 258
rect -272 105 -243 303
rect -525 23 -160 29
rect -525 -11 -480 23
rect -192 -11 -160 23
rect -525 -18 -160 -11
<< comment >>
rect -499 807 -1 808
rect -629 5 -526 6
rect -525 5 -160 6
rect -159 5 8 6
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_0
timestamp 1615245166
transform 1 0 -390 0 1 180
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_1
timestamp 1615245166
transform 1 0 -302 0 1 180
box -73 -116 73 116
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_0
timestamp 1615311486
transform 1 0 -390 0 1 627
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_1
timestamp 1615311486
transform 1 0 -302 0 1 627
box -109 -152 109 152
<< labels >>
rlabel metal1 -525 329 -453 357 1 A
rlabel metal1 -525 403 -300 431 1 B
rlabel nwell -463 788 -223 822 1 vdd
rlabel metal1 -456 -11 -216 23 1 vss
<< end >>
