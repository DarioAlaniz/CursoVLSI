magic
tech sky130A
magscale 1 2
timestamp 1614812053
<< error_p >>
rect -29 -161 29 -155
rect -29 -195 -17 -161
rect -29 -201 29 -195
<< nwell >>
rect -211 -334 211 334
<< pmos >>
rect -15 -114 15 186
<< pdiff >>
rect -73 174 -15 186
rect -73 -102 -61 174
rect -27 -102 -15 174
rect -73 -114 -15 -102
rect 15 174 73 186
rect 15 -102 27 174
rect 61 -102 73 174
rect 15 -114 73 -102
<< pdiffc >>
rect -61 -102 -27 174
rect 27 -102 61 174
<< nsubdiff >>
rect -175 264 -79 298
rect 79 264 175 298
rect -175 201 -141 264
rect 141 201 175 264
rect -175 -264 -141 -201
rect 141 -264 175 -201
rect -175 -298 175 -264
<< nsubdiffcont >>
rect -79 264 79 298
rect -175 -201 -141 201
rect 141 -201 175 201
<< poly >>
rect -15 186 15 212
rect -15 -145 15 -114
rect -33 -161 33 -145
rect -33 -195 -17 -161
rect 17 -195 33 -161
rect -33 -211 33 -195
<< polycont >>
rect -17 -195 17 -161
<< locali >>
rect -175 264 -79 298
rect 79 264 175 298
rect -175 201 -141 264
rect 141 201 175 264
rect -61 174 -27 190
rect -61 -118 -27 -102
rect 27 174 61 190
rect 27 -118 61 -102
rect -33 -195 -17 -161
rect 17 -195 33 -161
rect -175 -264 -141 -201
rect 141 -264 175 -201
rect -175 -298 175 -264
<< viali >>
rect -61 -102 -27 174
rect 27 -102 61 174
rect -17 -195 17 -161
<< metal1 >>
rect -67 174 -21 186
rect -67 -102 -61 174
rect -27 -102 -21 174
rect -67 -114 -21 -102
rect 21 174 67 186
rect 21 -102 27 174
rect 61 -102 67 174
rect 21 -114 67 -102
rect -29 -161 29 -155
rect -29 -195 -17 -161
rect 17 -195 29 -161
rect -29 -201 29 -195
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -158 -281 158 281
string parameters w 1.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
