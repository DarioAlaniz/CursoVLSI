magic
tech sky130A
magscale 1 2
timestamp 1615245166
<< error_p >>
rect -61 58 -27 64
rect -89 42 0 58
rect -89 30 1 42
rect -67 -12 -39 30
rect -27 -12 1 30
rect -67 -30 1 -12
rect -67 -42 -21 -30
rect -61 -46 -27 -42
<< nmos >>
rect -15 -42 15 60
<< ndiff >>
rect -73 -42 -15 60
rect 15 30 73 60
rect 15 -30 27 30
rect 61 -30 73 30
rect 15 -42 73 -30
<< ndiffc >>
rect 27 -30 61 30
<< poly >>
rect -15 60 15 86
rect -15 -68 15 -42
<< locali >>
rect -61 30 -27 46
rect 27 30 61 46
rect -61 -46 -27 -30
rect 27 -46 61 -30
<< viali >>
rect 27 -30 61 30
<< metal1 >>
rect -67 30 -21 42
rect -67 -30 -61 30
rect -27 -30 -21 30
rect -67 -42 -21 -30
rect 21 30 67 42
rect 21 -30 27 30
rect 61 -30 67 30
rect 21 -42 67 -30
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 0.420 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
